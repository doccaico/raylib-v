module math

#flag -I @VMODROOT/include

#include "raymath.h"
