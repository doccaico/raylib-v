module raymath

#flag -I @VMODROOT/include

#include "raymath.h"
