module gui

#flag -I @VMODROOT/include

#define RAYGUI_IMPLEMENTATION
#include "raygui.h"
